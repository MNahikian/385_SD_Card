// DE2_115_SD_CARD_NIOS.v

// Generated using ACDS version 14.1 186 at 2016.05.31.19:11:49

`timescale 1 ps / 1 ps
module DE2_115_SD_CARD_NIOS (
		input  wire        altpll_areset_conduit_export,                                    //               altpll_areset_conduit.export
		output wire        altpll_c1_clk,                                                   //                           altpll_c1.clk
		output wire        altpll_c3_clk,                                                   //                           altpll_c3.clk
		output wire        altpll_locked_conduit_export,                                    //               altpll_locked_conduit.export
		output wire        altpll_phasedone_conduit_export,                                 //            altpll_phasedone_conduit.export
		output wire        c0_out_clk_clk,                                                  //                          c0_out_clk.clk
		output wire        c2_out_clk_clk,                                                  //                          c2_out_clk.clk
		input  wire        clk_50_clk_in_clk,                                               //                       clk_50_clk_in.clk
		output wire        epp_i2c_scl_external_connection_export,                          //     epp_i2c_scl_external_connection.export
		inout  wire        epp_i2c_sda_external_connection_export,                          //     epp_i2c_sda_external_connection.export
		output wire        i2c_scl_external_connection_export,                              //         i2c_scl_external_connection.export
		inout  wire        i2c_sda_external_connection_export,                              //         i2c_sda_external_connection.export
		input  wire        ir_external_connection_export,                                   //              ir_external_connection.export
		input  wire [3:0]  key_external_connection_export,                                  //             key_external_connection.export
		output wire        lcd_external_RS,                                                 //                        lcd_external.RS
		output wire        lcd_external_RW,                                                 //                                    .RW
		inout  wire [7:0]  lcd_external_data,                                               //                                    .data
		output wire        lcd_external_E,                                                  //                                    .E
		output wire [8:0]  ledg_external_connection_export,                                 //            ledg_external_connection.export
		output wire [17:0] ledr_external_connection_export,                                 //            ledr_external_connection.export
		input  wire        reset_reset_n,                                                   //                               reset.reset_n
		input  wire        rs232_external_connection_rxd,                                   //           rs232_external_connection.rxd
		output wire        rs232_external_connection_txd,                                   //                                    .txd
		input  wire        rs232_external_connection_cts_n,                                 //                                    .cts_n
		output wire        rs232_external_connection_rts_n,                                 //                                    .rts_n
		output wire        sd_clk_external_connection_export,                               //          sd_clk_external_connection.export
		inout  wire        sd_cmd_external_connection_export,                               //          sd_cmd_external_connection.export
		inout  wire [3:0]  sd_dat_external_connection_export,                               //          sd_dat_external_connection.export
		input  wire        sd_wp_n_external_connection_export,                              //         sd_wp_n_external_connection.export
		output wire [63:0] seg7_conduit_end_export,                                         //                    seg7_conduit_end.export
		input  wire        sma_in_external_connection_export,                               //          sma_in_external_connection.export
		output wire        sma_out_external_connection_export,                              //         sma_out_external_connection.export
		input  wire [17:0] sw_external_connection_export,                                   //              sw_external_connection.export
		output wire [15:0] to_hw_port_export,                                               //                          to_hw_port.export
		output wire [1:0]  to_hw_sig_export,                                                //                           to_hw_sig.export
		input  wire [1:0]  to_sw_sig_export,                                                //                           to_sw_sig.export
		output wire [22:0] tri_state_bridge_flash_bridge_0_out_address_to_the_cfi_flash,    // tri_state_bridge_flash_bridge_0_out.address_to_the_cfi_flash
		inout  wire [7:0]  tri_state_bridge_flash_bridge_0_out_tri_state_bridge_flash_data, //                                    .tri_state_bridge_flash_data
		output wire [0:0]  tri_state_bridge_flash_bridge_0_out_write_n_to_the_cfi_flash,    //                                    .write_n_to_the_cfi_flash
		output wire [0:0]  tri_state_bridge_flash_bridge_0_out_select_n_to_the_cfi_flash,   //                                    .select_n_to_the_cfi_flash
		output wire [0:0]  tri_state_bridge_flash_bridge_0_out_read_n_to_the_cfi_flash      //                                    .read_n_to_the_cfi_flash
	);

	wire         cpu_jtag_debug_module_reset_reset;                                        // cpu:jtag_debug_module_resetrequest -> [epp_i2c_scl:reset_n, mm_interconnect_1:epp_i2c_scl_reset_reset_bridge_in_reset_reset, rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         tri_state_flash_bridge_pinsharer_0_tcm_request;                           // tri_state_flash_bridge_pinSharer_0:request -> tri_state_bridge_flash_bridge_0:request
	wire   [0:0] tri_state_flash_bridge_pinsharer_0_tcm_read_n_to_the_cfi_flash_out;       // tri_state_flash_bridge_pinSharer_0:read_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_read_n_to_the_cfi_flash
	wire  [22:0] tri_state_flash_bridge_pinsharer_0_tcm_address_to_the_cfi_flash_out;      // tri_state_flash_bridge_pinSharer_0:address_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_address_to_the_cfi_flash
	wire         tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_outen; // tri_state_flash_bridge_pinSharer_0:tri_state_bridge_flash_data_outen -> tri_state_bridge_flash_bridge_0:tcs_tri_state_bridge_flash_data_outen
	wire   [0:0] tri_state_flash_bridge_pinsharer_0_tcm_write_n_to_the_cfi_flash_out;      // tri_state_flash_bridge_pinSharer_0:write_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_write_n_to_the_cfi_flash
	wire   [7:0] tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_in;    // tri_state_bridge_flash_bridge_0:tcs_tri_state_bridge_flash_data_in -> tri_state_flash_bridge_pinSharer_0:tri_state_bridge_flash_data_in
	wire         tri_state_flash_bridge_pinsharer_0_tcm_grant;                             // tri_state_bridge_flash_bridge_0:grant -> tri_state_flash_bridge_pinSharer_0:grant
	wire   [7:0] tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_out;   // tri_state_flash_bridge_pinSharer_0:tri_state_bridge_flash_data -> tri_state_bridge_flash_bridge_0:tcs_tri_state_bridge_flash_data
	wire   [0:0] tri_state_flash_bridge_pinsharer_0_tcm_select_n_to_the_cfi_flash_out;     // tri_state_flash_bridge_pinSharer_0:select_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_select_n_to_the_cfi_flash
	wire         cfi_flash_tcm_data_outen;                                                 // cfi_flash:tcm_data_outen -> tri_state_flash_bridge_pinSharer_0:tcs0_data_outen
	wire         cfi_flash_tcm_request;                                                    // cfi_flash:tcm_request -> tri_state_flash_bridge_pinSharer_0:tcs0_request
	wire         cfi_flash_tcm_write_n_out;                                                // cfi_flash:tcm_write_n_out -> tri_state_flash_bridge_pinSharer_0:tcs0_write_n_out
	wire         cfi_flash_tcm_read_n_out;                                                 // cfi_flash:tcm_read_n_out -> tri_state_flash_bridge_pinSharer_0:tcs0_read_n_out
	wire         cfi_flash_tcm_grant;                                                      // tri_state_flash_bridge_pinSharer_0:tcs0_grant -> cfi_flash:tcm_grant
	wire         cfi_flash_tcm_chipselect_n_out;                                           // cfi_flash:tcm_chipselect_n_out -> tri_state_flash_bridge_pinSharer_0:tcs0_chipselect_n_out
	wire  [22:0] cfi_flash_tcm_address_out;                                                // cfi_flash:tcm_address_out -> tri_state_flash_bridge_pinSharer_0:tcs0_address_out
	wire   [7:0] cfi_flash_tcm_data_out;                                                   // cfi_flash:tcm_data_out -> tri_state_flash_bridge_pinSharer_0:tcs0_data_out
	wire   [7:0] cfi_flash_tcm_data_in;                                                    // tri_state_flash_bridge_pinSharer_0:tcs0_data_in -> cfi_flash:tcm_data_in
	wire  [31:0] cpu_data_master_readdata;                                                 // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                              // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                              // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [25:0] cpu_data_master_address;                                                  // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                               // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                     // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                                            // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                                    // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                                // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                          // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                       // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [25:0] cpu_instruction_master_address;                                           // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                              // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                                     // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                   // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                         // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;                      // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;                      // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                          // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                             // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;                       // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                            // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;                        // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_readdata;                              // altpll:readdata -> mm_interconnect_0:altpll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_pll_slave_address;                               // mm_interconnect_0:altpll_pll_slave_address -> altpll:address
	wire         mm_interconnect_0_altpll_pll_slave_read;                                  // mm_interconnect_0:altpll_pll_slave_read -> altpll:read
	wire         mm_interconnect_0_altpll_pll_slave_write;                                 // mm_interconnect_0:altpll_pll_slave_write -> altpll:write
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_writedata;                             // mm_interconnect_0:altpll_pll_slave_writedata -> altpll:writedata
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_readdata;                          // clock_crossing_io:s0_readdata -> mm_interconnect_0:clock_crossing_io_s0_readdata
	wire         mm_interconnect_0_clock_crossing_io_s0_waitrequest;                       // clock_crossing_io:s0_waitrequest -> mm_interconnect_0:clock_crossing_io_s0_waitrequest
	wire         mm_interconnect_0_clock_crossing_io_s0_debugaccess;                       // mm_interconnect_0:clock_crossing_io_s0_debugaccess -> clock_crossing_io:s0_debugaccess
	wire   [8:0] mm_interconnect_0_clock_crossing_io_s0_address;                           // mm_interconnect_0:clock_crossing_io_s0_address -> clock_crossing_io:s0_address
	wire         mm_interconnect_0_clock_crossing_io_s0_read;                              // mm_interconnect_0:clock_crossing_io_s0_read -> clock_crossing_io:s0_read
	wire   [3:0] mm_interconnect_0_clock_crossing_io_s0_byteenable;                        // mm_interconnect_0:clock_crossing_io_s0_byteenable -> clock_crossing_io:s0_byteenable
	wire         mm_interconnect_0_clock_crossing_io_s0_readdatavalid;                     // clock_crossing_io:s0_readdatavalid -> mm_interconnect_0:clock_crossing_io_s0_readdatavalid
	wire         mm_interconnect_0_clock_crossing_io_s0_write;                             // mm_interconnect_0:clock_crossing_io_s0_write -> clock_crossing_io:s0_write
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_writedata;                         // mm_interconnect_0:clock_crossing_io_s0_writedata -> clock_crossing_io:s0_writedata
	wire   [0:0] mm_interconnect_0_clock_crossing_io_s0_burstcount;                        // mm_interconnect_0:clock_crossing_io_s0_burstcount -> clock_crossing_io:s0_burstcount
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;                           // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;                             // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_s1_address;                              // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;                           // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                                // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;                            // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                                // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire  [31:0] mm_interconnect_0_sma_in_s1_readdata;                                     // sma_in:readdata -> mm_interconnect_0:sma_in_s1_readdata
	wire   [1:0] mm_interconnect_0_sma_in_s1_address;                                      // mm_interconnect_0:sma_in_s1_address -> sma_in:address
	wire         mm_interconnect_0_sma_out_s1_chipselect;                                  // mm_interconnect_0:sma_out_s1_chipselect -> sma_out:chipselect
	wire  [31:0] mm_interconnect_0_sma_out_s1_readdata;                                    // sma_out:readdata -> mm_interconnect_0:sma_out_s1_readdata
	wire   [1:0] mm_interconnect_0_sma_out_s1_address;                                     // mm_interconnect_0:sma_out_s1_address -> sma_out:address
	wire         mm_interconnect_0_sma_out_s1_write;                                       // mm_interconnect_0:sma_out_s1_write -> sma_out:write_n
	wire  [31:0] mm_interconnect_0_sma_out_s1_writedata;                                   // mm_interconnect_0:sma_out_s1_writedata -> sma_out:writedata
	wire   [7:0] mm_interconnect_0_cfi_flash_uas_readdata;                                 // cfi_flash:uas_readdata -> mm_interconnect_0:cfi_flash_uas_readdata
	wire         mm_interconnect_0_cfi_flash_uas_waitrequest;                              // cfi_flash:uas_waitrequest -> mm_interconnect_0:cfi_flash_uas_waitrequest
	wire         mm_interconnect_0_cfi_flash_uas_debugaccess;                              // mm_interconnect_0:cfi_flash_uas_debugaccess -> cfi_flash:uas_debugaccess
	wire  [22:0] mm_interconnect_0_cfi_flash_uas_address;                                  // mm_interconnect_0:cfi_flash_uas_address -> cfi_flash:uas_address
	wire         mm_interconnect_0_cfi_flash_uas_read;                                     // mm_interconnect_0:cfi_flash_uas_read -> cfi_flash:uas_read
	wire   [0:0] mm_interconnect_0_cfi_flash_uas_byteenable;                               // mm_interconnect_0:cfi_flash_uas_byteenable -> cfi_flash:uas_byteenable
	wire         mm_interconnect_0_cfi_flash_uas_readdatavalid;                            // cfi_flash:uas_readdatavalid -> mm_interconnect_0:cfi_flash_uas_readdatavalid
	wire         mm_interconnect_0_cfi_flash_uas_lock;                                     // mm_interconnect_0:cfi_flash_uas_lock -> cfi_flash:uas_lock
	wire         mm_interconnect_0_cfi_flash_uas_write;                                    // mm_interconnect_0:cfi_flash_uas_write -> cfi_flash:uas_write
	wire   [7:0] mm_interconnect_0_cfi_flash_uas_writedata;                                // mm_interconnect_0:cfi_flash_uas_writedata -> cfi_flash:uas_writedata
	wire   [0:0] mm_interconnect_0_cfi_flash_uas_burstcount;                               // mm_interconnect_0:cfi_flash_uas_burstcount -> cfi_flash:uas_burstcount
	wire         clock_crossing_io_m0_waitrequest;                                         // mm_interconnect_1:clock_crossing_io_m0_waitrequest -> clock_crossing_io:m0_waitrequest
	wire  [31:0] clock_crossing_io_m0_readdata;                                            // mm_interconnect_1:clock_crossing_io_m0_readdata -> clock_crossing_io:m0_readdata
	wire         clock_crossing_io_m0_debugaccess;                                         // clock_crossing_io:m0_debugaccess -> mm_interconnect_1:clock_crossing_io_m0_debugaccess
	wire   [8:0] clock_crossing_io_m0_address;                                             // clock_crossing_io:m0_address -> mm_interconnect_1:clock_crossing_io_m0_address
	wire         clock_crossing_io_m0_read;                                                // clock_crossing_io:m0_read -> mm_interconnect_1:clock_crossing_io_m0_read
	wire   [3:0] clock_crossing_io_m0_byteenable;                                          // clock_crossing_io:m0_byteenable -> mm_interconnect_1:clock_crossing_io_m0_byteenable
	wire         clock_crossing_io_m0_readdatavalid;                                       // mm_interconnect_1:clock_crossing_io_m0_readdatavalid -> clock_crossing_io:m0_readdatavalid
	wire  [31:0] clock_crossing_io_m0_writedata;                                           // clock_crossing_io:m0_writedata -> mm_interconnect_1:clock_crossing_io_m0_writedata
	wire         clock_crossing_io_m0_write;                                               // clock_crossing_io:m0_write -> mm_interconnect_1:clock_crossing_io_m0_write
	wire   [0:0] clock_crossing_io_m0_burstcount;                                          // clock_crossing_io:m0_burstcount -> mm_interconnect_1:clock_crossing_io_m0_burstcount
	wire   [7:0] mm_interconnect_1_seg7_avalon_slave_readdata;                             // seg7:s_readdata -> mm_interconnect_1:seg7_avalon_slave_readdata
	wire   [2:0] mm_interconnect_1_seg7_avalon_slave_address;                              // mm_interconnect_1:seg7_avalon_slave_address -> seg7:s_address
	wire         mm_interconnect_1_seg7_avalon_slave_read;                                 // mm_interconnect_1:seg7_avalon_slave_read -> seg7:s_read
	wire         mm_interconnect_1_seg7_avalon_slave_write;                                // mm_interconnect_1:seg7_avalon_slave_write -> seg7:s_write
	wire   [7:0] mm_interconnect_1_seg7_avalon_slave_writedata;                            // mm_interconnect_1:seg7_avalon_slave_writedata -> seg7:s_writedata
	wire   [7:0] mm_interconnect_1_lcd_control_slave_readdata;                             // lcd:readdata -> mm_interconnect_1:lcd_control_slave_readdata
	wire   [1:0] mm_interconnect_1_lcd_control_slave_address;                              // mm_interconnect_1:lcd_control_slave_address -> lcd:address
	wire         mm_interconnect_1_lcd_control_slave_read;                                 // mm_interconnect_1:lcd_control_slave_read -> lcd:read
	wire         mm_interconnect_1_lcd_control_slave_begintransfer;                        // mm_interconnect_1:lcd_control_slave_begintransfer -> lcd:begintransfer
	wire         mm_interconnect_1_lcd_control_slave_write;                                // mm_interconnect_1:lcd_control_slave_write -> lcd:write
	wire   [7:0] mm_interconnect_1_lcd_control_slave_writedata;                            // mm_interconnect_1:lcd_control_slave_writedata -> lcd:writedata
	wire         mm_interconnect_1_key_s1_chipselect;                                      // mm_interconnect_1:key_s1_chipselect -> key:chipselect
	wire  [31:0] mm_interconnect_1_key_s1_readdata;                                        // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire   [1:0] mm_interconnect_1_key_s1_address;                                         // mm_interconnect_1:key_s1_address -> key:address
	wire         mm_interconnect_1_key_s1_write;                                           // mm_interconnect_1:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_1_key_s1_writedata;                                       // mm_interconnect_1:key_s1_writedata -> key:writedata
	wire         mm_interconnect_1_sd_clk_s1_chipselect;                                   // mm_interconnect_1:sd_clk_s1_chipselect -> sd_clk:chipselect
	wire  [31:0] mm_interconnect_1_sd_clk_s1_readdata;                                     // sd_clk:readdata -> mm_interconnect_1:sd_clk_s1_readdata
	wire   [1:0] mm_interconnect_1_sd_clk_s1_address;                                      // mm_interconnect_1:sd_clk_s1_address -> sd_clk:address
	wire         mm_interconnect_1_sd_clk_s1_write;                                        // mm_interconnect_1:sd_clk_s1_write -> sd_clk:write_n
	wire  [31:0] mm_interconnect_1_sd_clk_s1_writedata;                                    // mm_interconnect_1:sd_clk_s1_writedata -> sd_clk:writedata
	wire         mm_interconnect_1_sd_cmd_s1_chipselect;                                   // mm_interconnect_1:sd_cmd_s1_chipselect -> sd_cmd:chipselect
	wire  [31:0] mm_interconnect_1_sd_cmd_s1_readdata;                                     // sd_cmd:readdata -> mm_interconnect_1:sd_cmd_s1_readdata
	wire   [1:0] mm_interconnect_1_sd_cmd_s1_address;                                      // mm_interconnect_1:sd_cmd_s1_address -> sd_cmd:address
	wire         mm_interconnect_1_sd_cmd_s1_write;                                        // mm_interconnect_1:sd_cmd_s1_write -> sd_cmd:write_n
	wire  [31:0] mm_interconnect_1_sd_cmd_s1_writedata;                                    // mm_interconnect_1:sd_cmd_s1_writedata -> sd_cmd:writedata
	wire         mm_interconnect_1_sd_dat_s1_chipselect;                                   // mm_interconnect_1:sd_dat_s1_chipselect -> sd_dat:chipselect
	wire  [31:0] mm_interconnect_1_sd_dat_s1_readdata;                                     // sd_dat:readdata -> mm_interconnect_1:sd_dat_s1_readdata
	wire   [1:0] mm_interconnect_1_sd_dat_s1_address;                                      // mm_interconnect_1:sd_dat_s1_address -> sd_dat:address
	wire         mm_interconnect_1_sd_dat_s1_write;                                        // mm_interconnect_1:sd_dat_s1_write -> sd_dat:write_n
	wire  [31:0] mm_interconnect_1_sd_dat_s1_writedata;                                    // mm_interconnect_1:sd_dat_s1_writedata -> sd_dat:writedata
	wire  [31:0] mm_interconnect_1_sd_wp_n_s1_readdata;                                    // sd_wp_n:readdata -> mm_interconnect_1:sd_wp_n_s1_readdata
	wire   [1:0] mm_interconnect_1_sd_wp_n_s1_address;                                     // mm_interconnect_1:sd_wp_n_s1_address -> sd_wp_n:address
	wire         mm_interconnect_1_epp_i2c_scl_s1_chipselect;                              // mm_interconnect_1:epp_i2c_scl_s1_chipselect -> epp_i2c_scl:chipselect
	wire  [31:0] mm_interconnect_1_epp_i2c_scl_s1_readdata;                                // epp_i2c_scl:readdata -> mm_interconnect_1:epp_i2c_scl_s1_readdata
	wire   [1:0] mm_interconnect_1_epp_i2c_scl_s1_address;                                 // mm_interconnect_1:epp_i2c_scl_s1_address -> epp_i2c_scl:address
	wire         mm_interconnect_1_epp_i2c_scl_s1_write;                                   // mm_interconnect_1:epp_i2c_scl_s1_write -> epp_i2c_scl:write_n
	wire  [31:0] mm_interconnect_1_epp_i2c_scl_s1_writedata;                               // mm_interconnect_1:epp_i2c_scl_s1_writedata -> epp_i2c_scl:writedata
	wire         mm_interconnect_1_epp_i2c_sda_s1_chipselect;                              // mm_interconnect_1:epp_i2c_sda_s1_chipselect -> epp_i2c_sda:chipselect
	wire  [31:0] mm_interconnect_1_epp_i2c_sda_s1_readdata;                                // epp_i2c_sda:readdata -> mm_interconnect_1:epp_i2c_sda_s1_readdata
	wire   [1:0] mm_interconnect_1_epp_i2c_sda_s1_address;                                 // mm_interconnect_1:epp_i2c_sda_s1_address -> epp_i2c_sda:address
	wire         mm_interconnect_1_epp_i2c_sda_s1_write;                                   // mm_interconnect_1:epp_i2c_sda_s1_write -> epp_i2c_sda:write_n
	wire  [31:0] mm_interconnect_1_epp_i2c_sda_s1_writedata;                               // mm_interconnect_1:epp_i2c_sda_s1_writedata -> epp_i2c_sda:writedata
	wire         mm_interconnect_1_sw_s1_chipselect;                                       // mm_interconnect_1:sw_s1_chipselect -> sw:chipselect
	wire  [31:0] mm_interconnect_1_sw_s1_readdata;                                         // sw:readdata -> mm_interconnect_1:sw_s1_readdata
	wire   [1:0] mm_interconnect_1_sw_s1_address;                                          // mm_interconnect_1:sw_s1_address -> sw:address
	wire         mm_interconnect_1_sw_s1_write;                                            // mm_interconnect_1:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_1_sw_s1_writedata;                                        // mm_interconnect_1:sw_s1_writedata -> sw:writedata
	wire         mm_interconnect_1_i2c_scl_s1_chipselect;                                  // mm_interconnect_1:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	wire  [31:0] mm_interconnect_1_i2c_scl_s1_readdata;                                    // i2c_scl:readdata -> mm_interconnect_1:i2c_scl_s1_readdata
	wire   [1:0] mm_interconnect_1_i2c_scl_s1_address;                                     // mm_interconnect_1:i2c_scl_s1_address -> i2c_scl:address
	wire         mm_interconnect_1_i2c_scl_s1_write;                                       // mm_interconnect_1:i2c_scl_s1_write -> i2c_scl:write_n
	wire  [31:0] mm_interconnect_1_i2c_scl_s1_writedata;                                   // mm_interconnect_1:i2c_scl_s1_writedata -> i2c_scl:writedata
	wire         mm_interconnect_1_i2c_sda_s1_chipselect;                                  // mm_interconnect_1:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	wire  [31:0] mm_interconnect_1_i2c_sda_s1_readdata;                                    // i2c_sda:readdata -> mm_interconnect_1:i2c_sda_s1_readdata
	wire   [1:0] mm_interconnect_1_i2c_sda_s1_address;                                     // mm_interconnect_1:i2c_sda_s1_address -> i2c_sda:address
	wire         mm_interconnect_1_i2c_sda_s1_write;                                       // mm_interconnect_1:i2c_sda_s1_write -> i2c_sda:write_n
	wire  [31:0] mm_interconnect_1_i2c_sda_s1_writedata;                                   // mm_interconnect_1:i2c_sda_s1_writedata -> i2c_sda:writedata
	wire         mm_interconnect_1_timer_s1_chipselect;                                    // mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_1_timer_s1_readdata;                                      // timer:readdata -> mm_interconnect_1:timer_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_s1_address;                                       // mm_interconnect_1:timer_s1_address -> timer:address
	wire         mm_interconnect_1_timer_s1_write;                                         // mm_interconnect_1:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_1_timer_s1_writedata;                                     // mm_interconnect_1:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_1_ledg_s1_chipselect;                                     // mm_interconnect_1:ledg_s1_chipselect -> ledg:chipselect
	wire  [31:0] mm_interconnect_1_ledg_s1_readdata;                                       // ledg:readdata -> mm_interconnect_1:ledg_s1_readdata
	wire   [1:0] mm_interconnect_1_ledg_s1_address;                                        // mm_interconnect_1:ledg_s1_address -> ledg:address
	wire         mm_interconnect_1_ledg_s1_write;                                          // mm_interconnect_1:ledg_s1_write -> ledg:write_n
	wire  [31:0] mm_interconnect_1_ledg_s1_writedata;                                      // mm_interconnect_1:ledg_s1_writedata -> ledg:writedata
	wire         mm_interconnect_1_ledr_s1_chipselect;                                     // mm_interconnect_1:ledr_s1_chipselect -> ledr:chipselect
	wire  [31:0] mm_interconnect_1_ledr_s1_readdata;                                       // ledr:readdata -> mm_interconnect_1:ledr_s1_readdata
	wire   [1:0] mm_interconnect_1_ledr_s1_address;                                        // mm_interconnect_1:ledr_s1_address -> ledr:address
	wire         mm_interconnect_1_ledr_s1_write;                                          // mm_interconnect_1:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_1_ledr_s1_writedata;                                      // mm_interconnect_1:ledr_s1_writedata -> ledr:writedata
	wire  [31:0] mm_interconnect_1_ir_s1_readdata;                                         // ir:readdata -> mm_interconnect_1:ir_s1_readdata
	wire   [1:0] mm_interconnect_1_ir_s1_address;                                          // mm_interconnect_1:ir_s1_address -> ir:address
	wire         mm_interconnect_1_rs232_s1_chipselect;                                    // mm_interconnect_1:rs232_s1_chipselect -> rs232:chipselect
	wire  [15:0] mm_interconnect_1_rs232_s1_readdata;                                      // rs232:readdata -> mm_interconnect_1:rs232_s1_readdata
	wire   [2:0] mm_interconnect_1_rs232_s1_address;                                       // mm_interconnect_1:rs232_s1_address -> rs232:address
	wire         mm_interconnect_1_rs232_s1_read;                                          // mm_interconnect_1:rs232_s1_read -> rs232:read_n
	wire         mm_interconnect_1_rs232_s1_begintransfer;                                 // mm_interconnect_1:rs232_s1_begintransfer -> rs232:begintransfer
	wire         mm_interconnect_1_rs232_s1_write;                                         // mm_interconnect_1:rs232_s1_write -> rs232:write_n
	wire  [15:0] mm_interconnect_1_rs232_s1_writedata;                                     // mm_interconnect_1:rs232_s1_writedata -> rs232:writedata
	wire  [31:0] mm_interconnect_1_to_sw_sig_s1_readdata;                                  // to_sw_sig:readdata -> mm_interconnect_1:to_sw_sig_s1_readdata
	wire   [1:0] mm_interconnect_1_to_sw_sig_s1_address;                                   // mm_interconnect_1:to_sw_sig_s1_address -> to_sw_sig:address
	wire         mm_interconnect_1_to_hw_sig_s1_chipselect;                                // mm_interconnect_1:to_hw_sig_s1_chipselect -> to_hw_sig:chipselect
	wire  [31:0] mm_interconnect_1_to_hw_sig_s1_readdata;                                  // to_hw_sig:readdata -> mm_interconnect_1:to_hw_sig_s1_readdata
	wire   [1:0] mm_interconnect_1_to_hw_sig_s1_address;                                   // mm_interconnect_1:to_hw_sig_s1_address -> to_hw_sig:address
	wire         mm_interconnect_1_to_hw_sig_s1_write;                                     // mm_interconnect_1:to_hw_sig_s1_write -> to_hw_sig:write_n
	wire  [31:0] mm_interconnect_1_to_hw_sig_s1_writedata;                                 // mm_interconnect_1:to_hw_sig_s1_writedata -> to_hw_sig:writedata
	wire         mm_interconnect_1_to_hw_port_s1_chipselect;                               // mm_interconnect_1:to_hw_port_s1_chipselect -> to_hw_port:chipselect
	wire  [31:0] mm_interconnect_1_to_hw_port_s1_readdata;                                 // to_hw_port:readdata -> mm_interconnect_1:to_hw_port_s1_readdata
	wire   [1:0] mm_interconnect_1_to_hw_port_s1_address;                                  // mm_interconnect_1:to_hw_port_s1_address -> to_hw_port:address
	wire         mm_interconnect_1_to_hw_port_s1_write;                                    // mm_interconnect_1:to_hw_port_s1_write -> to_hw_port:write_n
	wire  [31:0] mm_interconnect_1_to_hw_port_s1_writedata;                                // mm_interconnect_1:to_hw_port_s1_writedata -> to_hw_port:writedata
	wire         irq_mapper_receiver0_irq;                                                 // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                 // key:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                 // sw:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                 // rs232:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                 // timer:irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_d_irq_irq;                                                            // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                                           // rst_controller:reset_out -> [altpll:reset, mm_interconnect_0:altpll_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                       // rst_controller_001:reset_out -> [cfi_flash:reset_reset, clock_crossing_io:s0_reset, cpu:reset_n, epp_i2c_sda:reset_n, i2c_scl:reset_n, i2c_sda:reset_n, irq_mapper:reset, jtag_uart:rst_n, key:reset_n, lcd:reset_n, ledg:reset_n, ledr:reset_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:seg7_clock_sink_reset_reset_bridge_in_reset_reset, rs232:reset_n, rst_translator:in_reset, sd_clk:reset_n, sd_cmd:reset_n, sd_dat:reset_n, sd_wp_n:reset_n, seg7:s_reset, sma_in:reset_n, sma_out:reset_n, sw:reset_n, timer:reset_n, to_hw_port:reset_n, to_hw_sig:reset_n, to_sw_sig:reset_n, tri_state_bridge_flash_bridge_0:reset, tri_state_flash_bridge_pinSharer_0:reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                                   // rst_controller_001:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                                       // rst_controller_002:reset_out -> [clock_crossing_io:m0_reset, mm_interconnect_1:clock_crossing_io_m0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_003_reset_out_reset;                                       // rst_controller_003:reset_out -> [ir:reset_n, mm_interconnect_0:onchip_memory2_reset1_reset_bridge_in_reset_reset, mm_interconnect_1:ir_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_translator_001:in_reset]
	wire         rst_controller_003_reset_out_reset_req;                                   // rst_controller_003:reset_req -> [onchip_memory2:reset_req, rst_translator_001:reset_req_in]

	DE2_115_SD_CARD_NIOS_altpll altpll (
		.clk       (clk_50_clk_in_clk),                            //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),               // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_pll_slave_writedata), //                      .writedata
		.c0        (c0_out_clk_clk),                               //                    c0.clk
		.c1        (altpll_c1_clk),                                //                    c1.clk
		.c2        (c2_out_clk_clk),                               //                    c2.clk
		.c3        (altpll_c3_clk),                                //                    c3.clk
		.areset    (altpll_areset_conduit_export),                 //        areset_conduit.export
		.locked    (altpll_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (altpll_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	DE2_115_SD_CARD_NIOS_cfi_flash #(
		.TCM_ADDRESS_W                  (23),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (0),
		.TCM_WRITE_WAIT                 (0),
		.TCM_SETUP_WAIT                 (0),
		.TCM_DATA_HOLD                  (0),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) cfi_flash (
		.clk_clk              (c0_out_clk_clk),                                //   clk.clk
		.reset_reset          (rst_controller_001_reset_out_reset),            // reset.reset
		.uas_address          (mm_interconnect_0_cfi_flash_uas_address),       //   uas.address
		.uas_burstcount       (mm_interconnect_0_cfi_flash_uas_burstcount),    //      .burstcount
		.uas_read             (mm_interconnect_0_cfi_flash_uas_read),          //      .read
		.uas_write            (mm_interconnect_0_cfi_flash_uas_write),         //      .write
		.uas_waitrequest      (mm_interconnect_0_cfi_flash_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (mm_interconnect_0_cfi_flash_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable       (mm_interconnect_0_cfi_flash_uas_byteenable),    //      .byteenable
		.uas_readdata         (mm_interconnect_0_cfi_flash_uas_readdata),      //      .readdata
		.uas_writedata        (mm_interconnect_0_cfi_flash_uas_writedata),     //      .writedata
		.uas_lock             (mm_interconnect_0_cfi_flash_uas_lock),          //      .lock
		.uas_debugaccess      (mm_interconnect_0_cfi_flash_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (cfi_flash_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_read_n_out       (cfi_flash_tcm_read_n_out),                      //      .read_n_out
		.tcm_chipselect_n_out (cfi_flash_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_request          (cfi_flash_tcm_request),                         //      .request
		.tcm_grant            (cfi_flash_tcm_grant),                           //      .grant
		.tcm_address_out      (cfi_flash_tcm_address_out),                     //      .address_out
		.tcm_data_out         (cfi_flash_tcm_data_out),                        //      .data_out
		.tcm_data_outen       (cfi_flash_tcm_data_outen),                      //      .data_outen
		.tcm_data_in          (cfi_flash_tcm_data_in)                          //      .data_in
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (9),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (256),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_io (
		.m0_clk           (c2_out_clk_clk),                                       //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                   // m0_reset.reset
		.s0_clk           (c0_out_clk_clk),                                       //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                   // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_clock_crossing_io_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_clock_crossing_io_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_clock_crossing_io_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_clock_crossing_io_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_clock_crossing_io_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_clock_crossing_io_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_clock_crossing_io_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_clock_crossing_io_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_clock_crossing_io_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_clock_crossing_io_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_io_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_io_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_io_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_io_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_io_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_io_m0_address),                         //         .address
		.m0_write         (clock_crossing_io_m0_write),                           //         .write
		.m0_read          (clock_crossing_io_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_io_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_io_m0_debugaccess)                      //         .debugaccess
	);

	DE2_115_SD_CARD_NIOS_cpu cpu (
		.clk                                   (c0_out_clk_clk),                                      //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	DE2_115_SD_CARD_NIOS_epp_i2c_scl epp_i2c_scl (
		.clk        (c0_out_clk_clk),                              //                 clk.clk
		.reset_n    (~cpu_jtag_debug_module_reset_reset),          //               reset.reset_n
		.address    (mm_interconnect_1_epp_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_epp_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_epp_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_epp_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_epp_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (epp_i2c_scl_external_connection_export)       // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_epp_i2c_sda epp_i2c_sda (
		.clk        (c0_out_clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_epp_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_epp_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_epp_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_epp_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_epp_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (epp_i2c_sda_external_connection_export)       // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_epp_i2c_scl i2c_scl (
		.clk        (c0_out_clk_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (i2c_scl_external_connection_export)       // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_epp_i2c_sda i2c_sda (
		.clk        (c0_out_clk_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (i2c_sda_external_connection_export)       // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_ir ir (
		.clk      (c0_out_clk_clk),                      //                 clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_1_ir_s1_address),     //                  s1.address
		.readdata (mm_interconnect_1_ir_s1_readdata),    //                    .readdata
		.in_port  (ir_external_connection_export)        // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_jtag_uart jtag_uart (
		.clk            (c0_out_clk_clk),                                            //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	DE2_115_SD_CARD_NIOS_key key (
		.clk        (c0_out_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver1_irq)             //                 irq.irq
	);

	DE2_115_SD_CARD_NIOS_lcd lcd (
		.reset_n       (~rst_controller_001_reset_out_reset),               //         reset.reset_n
		.clk           (c0_out_clk_clk),                                    //           clk.clk
		.begintransfer (mm_interconnect_1_lcd_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_1_lcd_control_slave_read),          //              .read
		.write         (mm_interconnect_1_lcd_control_slave_write),         //              .write
		.readdata      (mm_interconnect_1_lcd_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_1_lcd_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_1_lcd_control_slave_address),       //              .address
		.LCD_RS        (lcd_external_RS),                                   //      external.export
		.LCD_RW        (lcd_external_RW),                                   //              .export
		.LCD_data      (lcd_external_data),                                 //              .export
		.LCD_E         (lcd_external_E)                                     //              .export
	);

	DE2_115_SD_CARD_NIOS_ledg ledg (
		.clk        (c0_out_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_1_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_external_connection_export)       // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_ledr ledr (
		.clk        (c0_out_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_1_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_external_connection_export)       // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_onchip_memory2 onchip_memory2 (
		.clk        (c0_out_clk_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_003_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_003_reset_out_reset_req)          //       .reset_req
	);

	DE2_115_SD_CARD_NIOS_rs232 rs232 (
		.clk           (c0_out_clk_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address       (mm_interconnect_1_rs232_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_1_rs232_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_1_rs232_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_1_rs232_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_1_rs232_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_1_rs232_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_1_rs232_s1_readdata),      //                    .readdata
		.dataavailable (),                                         //                    .dataavailable
		.readyfordata  (),                                         //                    .readyfordata
		.rxd           (rs232_external_connection_rxd),            // external_connection.export
		.txd           (rs232_external_connection_txd),            //                    .export
		.cts_n         (rs232_external_connection_cts_n),          //                    .export
		.rts_n         (rs232_external_connection_rts_n),          //                    .export
		.irq           (irq_mapper_receiver3_irq)                  //                 irq.irq
	);

	DE2_115_SD_CARD_NIOS_epp_i2c_scl sd_clk (
		.clk        (c0_out_clk_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sd_clk_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_clk_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_clk_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_clk_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_clk_s1_readdata),   //                    .readdata
		.out_port   (sd_clk_external_connection_export)       // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_epp_i2c_sda sd_cmd (
		.clk        (c0_out_clk_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sd_cmd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_cmd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_cmd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_cmd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_cmd_s1_readdata),   //                    .readdata
		.bidir_port (sd_cmd_external_connection_export)       // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_sd_dat sd_dat (
		.clk        (c0_out_clk_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sd_dat_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_dat_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_dat_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_dat_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_dat_s1_readdata),   //                    .readdata
		.bidir_port (sd_dat_external_connection_export)       // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_ir sd_wp_n (
		.clk      (c0_out_clk_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_1_sd_wp_n_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_sd_wp_n_s1_readdata), //                    .readdata
		.in_port  (sd_wp_n_external_connection_export)     // external_connection.export
	);

	SEG7_IF #(
		.SEG7_NUM       (8),
		.ADDR_WIDTH     (3),
		.DEFAULT_ACTIVE (1),
		.LOW_ACTIVE     (1)
	) seg7 (
		.s_address   (mm_interconnect_1_seg7_avalon_slave_address),   //     avalon_slave.address
		.s_read      (mm_interconnect_1_seg7_avalon_slave_read),      //                 .read
		.s_readdata  (mm_interconnect_1_seg7_avalon_slave_readdata),  //                 .readdata
		.s_write     (mm_interconnect_1_seg7_avalon_slave_write),     //                 .write
		.s_writedata (mm_interconnect_1_seg7_avalon_slave_writedata), //                 .writedata
		.SEG7        (seg7_conduit_end_export),                       //      conduit_end.export
		.s_clk       (c0_out_clk_clk),                                //       clock_sink.clk
		.s_reset     (rst_controller_001_reset_out_reset)             // clock_sink_reset.reset
	);

	DE2_115_SD_CARD_NIOS_ir sma_in (
		.clk      (c0_out_clk_clk),                       //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sma_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sma_in_s1_readdata), //                    .readdata
		.in_port  (sma_in_external_connection_export)     // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_epp_i2c_scl sma_out (
		.clk        (c0_out_clk_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_sma_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sma_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sma_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sma_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sma_out_s1_readdata),   //                    .readdata
		.out_port   (sma_out_external_connection_export)       // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_sw sw (
		.clk        (c0_out_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_sw_s1_address),     //                  s1.address
		.write_n    (~mm_interconnect_1_sw_s1_write),      //                    .write_n
		.writedata  (mm_interconnect_1_sw_s1_writedata),   //                    .writedata
		.chipselect (mm_interconnect_1_sw_s1_chipselect),  //                    .chipselect
		.readdata   (mm_interconnect_1_sw_s1_readdata),    //                    .readdata
		.in_port    (sw_external_connection_export),       // external_connection.export
		.irq        (irq_mapper_receiver2_irq)             //                 irq.irq
	);

	DE2_115_SD_CARD_NIOS_timer timer (
		.clk        (c0_out_clk_clk),                        //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_1_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)               //   irq.irq
	);

	DE2_115_SD_CARD_NIOS_to_hw_port to_hw_port (
		.clk        (c0_out_clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_1_to_hw_port_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_to_hw_port_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_to_hw_port_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_to_hw_port_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_to_hw_port_s1_readdata),   //                    .readdata
		.out_port   (to_hw_port_export)                           // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_to_hw_sig to_hw_sig (
		.clk        (c0_out_clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_1_to_hw_sig_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_to_hw_sig_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_to_hw_sig_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_to_hw_sig_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_to_hw_sig_s1_readdata),   //                    .readdata
		.out_port   (to_hw_sig_export)                           // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_to_sw_sig to_sw_sig (
		.clk      (c0_out_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_1_to_sw_sig_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_to_sw_sig_s1_readdata), //                    .readdata
		.in_port  (to_sw_sig_export)                         // external_connection.export
	);

	DE2_115_SD_CARD_NIOS_tri_state_bridge_flash_bridge_0 tri_state_bridge_flash_bridge_0 (
		.clk                                   (c0_out_clk_clk),                                                           //   clk.clk
		.reset                                 (rst_controller_001_reset_out_reset),                                       // reset.reset
		.request                               (tri_state_flash_bridge_pinsharer_0_tcm_request),                           //   tcs.request
		.grant                                 (tri_state_flash_bridge_pinsharer_0_tcm_grant),                             //      .grant
		.tcs_address_to_the_cfi_flash          (tri_state_flash_bridge_pinsharer_0_tcm_address_to_the_cfi_flash_out),      //      .address_to_the_cfi_flash_out
		.tcs_tri_state_bridge_flash_data       (tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_out),   //      .tri_state_bridge_flash_data_out
		.tcs_tri_state_bridge_flash_data_outen (tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_outen), //      .tri_state_bridge_flash_data_outen
		.tcs_tri_state_bridge_flash_data_in    (tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_in),    //      .tri_state_bridge_flash_data_in
		.tcs_write_n_to_the_cfi_flash          (tri_state_flash_bridge_pinsharer_0_tcm_write_n_to_the_cfi_flash_out),      //      .write_n_to_the_cfi_flash_out
		.tcs_select_n_to_the_cfi_flash         (tri_state_flash_bridge_pinsharer_0_tcm_select_n_to_the_cfi_flash_out),     //      .select_n_to_the_cfi_flash_out
		.tcs_read_n_to_the_cfi_flash           (tri_state_flash_bridge_pinsharer_0_tcm_read_n_to_the_cfi_flash_out),       //      .read_n_to_the_cfi_flash_out
		.address_to_the_cfi_flash              (tri_state_bridge_flash_bridge_0_out_address_to_the_cfi_flash),             //   out.address_to_the_cfi_flash
		.tri_state_bridge_flash_data           (tri_state_bridge_flash_bridge_0_out_tri_state_bridge_flash_data),          //      .tri_state_bridge_flash_data
		.write_n_to_the_cfi_flash              (tri_state_bridge_flash_bridge_0_out_write_n_to_the_cfi_flash),             //      .write_n_to_the_cfi_flash
		.select_n_to_the_cfi_flash             (tri_state_bridge_flash_bridge_0_out_select_n_to_the_cfi_flash),            //      .select_n_to_the_cfi_flash
		.read_n_to_the_cfi_flash               (tri_state_bridge_flash_bridge_0_out_read_n_to_the_cfi_flash)               //      .read_n_to_the_cfi_flash
	);

	DE2_115_SD_CARD_NIOS_tri_state_flash_bridge_pinSharer_0 tri_state_flash_bridge_pinsharer_0 (
		.clk_clk                           (c0_out_clk_clk),                                                           //   clk.clk
		.reset_reset                       (rst_controller_001_reset_out_reset),                                       // reset.reset
		.request                           (tri_state_flash_bridge_pinsharer_0_tcm_request),                           //   tcm.request
		.grant                             (tri_state_flash_bridge_pinsharer_0_tcm_grant),                             //      .grant
		.address_to_the_cfi_flash          (tri_state_flash_bridge_pinsharer_0_tcm_address_to_the_cfi_flash_out),      //      .address_to_the_cfi_flash_out
		.read_n_to_the_cfi_flash           (tri_state_flash_bridge_pinsharer_0_tcm_read_n_to_the_cfi_flash_out),       //      .read_n_to_the_cfi_flash_out
		.write_n_to_the_cfi_flash          (tri_state_flash_bridge_pinsharer_0_tcm_write_n_to_the_cfi_flash_out),      //      .write_n_to_the_cfi_flash_out
		.tri_state_bridge_flash_data       (tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_out),   //      .tri_state_bridge_flash_data_out
		.tri_state_bridge_flash_data_in    (tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_in),    //      .tri_state_bridge_flash_data_in
		.tri_state_bridge_flash_data_outen (tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_outen), //      .tri_state_bridge_flash_data_outen
		.select_n_to_the_cfi_flash         (tri_state_flash_bridge_pinsharer_0_tcm_select_n_to_the_cfi_flash_out),     //      .select_n_to_the_cfi_flash_out
		.tcs0_request                      (cfi_flash_tcm_request),                                                    //  tcs0.request
		.tcs0_grant                        (cfi_flash_tcm_grant),                                                      //      .grant
		.tcs0_address_out                  (cfi_flash_tcm_address_out),                                                //      .address_out
		.tcs0_read_n_out                   (cfi_flash_tcm_read_n_out),                                                 //      .read_n_out
		.tcs0_write_n_out                  (cfi_flash_tcm_write_n_out),                                                //      .write_n_out
		.tcs0_data_out                     (cfi_flash_tcm_data_out),                                                   //      .data_out
		.tcs0_data_in                      (cfi_flash_tcm_data_in),                                                    //      .data_in
		.tcs0_data_outen                   (cfi_flash_tcm_data_outen),                                                 //      .data_outen
		.tcs0_chipselect_n_out             (cfi_flash_tcm_chipselect_n_out)                                            //      .chipselect_n_out
	);

	DE2_115_SD_CARD_NIOS_mm_interconnect_0 mm_interconnect_0 (
		.altpll_c0_clk                                            (c0_out_clk_clk),                                            //                                          altpll_c0.clk
		.clk_50_clk_clk                                           (clk_50_clk_in_clk),                                         //                                         clk_50_clk.clk
		.altpll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // altpll_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_reset_n_reset_bridge_in_reset_reset                  (rst_controller_001_reset_out_reset),                        //                  cpu_reset_n_reset_bridge_in_reset.reset
		.onchip_memory2_reset1_reset_bridge_in_reset_reset        (rst_controller_003_reset_out_reset),                        //        onchip_memory2_reset1_reset_bridge_in_reset.reset
		.cpu_data_master_address                                  (cpu_data_master_address),                                   //                                    cpu_data_master.address
		.cpu_data_master_waitrequest                              (cpu_data_master_waitrequest),                               //                                                   .waitrequest
		.cpu_data_master_byteenable                               (cpu_data_master_byteenable),                                //                                                   .byteenable
		.cpu_data_master_read                                     (cpu_data_master_read),                                      //                                                   .read
		.cpu_data_master_readdata                                 (cpu_data_master_readdata),                                  //                                                   .readdata
		.cpu_data_master_readdatavalid                            (cpu_data_master_readdatavalid),                             //                                                   .readdatavalid
		.cpu_data_master_write                                    (cpu_data_master_write),                                     //                                                   .write
		.cpu_data_master_writedata                                (cpu_data_master_writedata),                                 //                                                   .writedata
		.cpu_data_master_debugaccess                              (cpu_data_master_debugaccess),                               //                                                   .debugaccess
		.cpu_instruction_master_address                           (cpu_instruction_master_address),                            //                             cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                       (cpu_instruction_master_waitrequest),                        //                                                   .waitrequest
		.cpu_instruction_master_read                              (cpu_instruction_master_read),                               //                                                   .read
		.cpu_instruction_master_readdata                          (cpu_instruction_master_readdata),                           //                                                   .readdata
		.cpu_instruction_master_readdatavalid                     (cpu_instruction_master_readdatavalid),                      //                                                   .readdatavalid
		.altpll_pll_slave_address                                 (mm_interconnect_0_altpll_pll_slave_address),                //                                   altpll_pll_slave.address
		.altpll_pll_slave_write                                   (mm_interconnect_0_altpll_pll_slave_write),                  //                                                   .write
		.altpll_pll_slave_read                                    (mm_interconnect_0_altpll_pll_slave_read),                   //                                                   .read
		.altpll_pll_slave_readdata                                (mm_interconnect_0_altpll_pll_slave_readdata),               //                                                   .readdata
		.altpll_pll_slave_writedata                               (mm_interconnect_0_altpll_pll_slave_writedata),              //                                                   .writedata
		.cfi_flash_uas_address                                    (mm_interconnect_0_cfi_flash_uas_address),                   //                                      cfi_flash_uas.address
		.cfi_flash_uas_write                                      (mm_interconnect_0_cfi_flash_uas_write),                     //                                                   .write
		.cfi_flash_uas_read                                       (mm_interconnect_0_cfi_flash_uas_read),                      //                                                   .read
		.cfi_flash_uas_readdata                                   (mm_interconnect_0_cfi_flash_uas_readdata),                  //                                                   .readdata
		.cfi_flash_uas_writedata                                  (mm_interconnect_0_cfi_flash_uas_writedata),                 //                                                   .writedata
		.cfi_flash_uas_burstcount                                 (mm_interconnect_0_cfi_flash_uas_burstcount),                //                                                   .burstcount
		.cfi_flash_uas_byteenable                                 (mm_interconnect_0_cfi_flash_uas_byteenable),                //                                                   .byteenable
		.cfi_flash_uas_readdatavalid                              (mm_interconnect_0_cfi_flash_uas_readdatavalid),             //                                                   .readdatavalid
		.cfi_flash_uas_waitrequest                                (mm_interconnect_0_cfi_flash_uas_waitrequest),               //                                                   .waitrequest
		.cfi_flash_uas_lock                                       (mm_interconnect_0_cfi_flash_uas_lock),                      //                                                   .lock
		.cfi_flash_uas_debugaccess                                (mm_interconnect_0_cfi_flash_uas_debugaccess),               //                                                   .debugaccess
		.clock_crossing_io_s0_address                             (mm_interconnect_0_clock_crossing_io_s0_address),            //                               clock_crossing_io_s0.address
		.clock_crossing_io_s0_write                               (mm_interconnect_0_clock_crossing_io_s0_write),              //                                                   .write
		.clock_crossing_io_s0_read                                (mm_interconnect_0_clock_crossing_io_s0_read),               //                                                   .read
		.clock_crossing_io_s0_readdata                            (mm_interconnect_0_clock_crossing_io_s0_readdata),           //                                                   .readdata
		.clock_crossing_io_s0_writedata                           (mm_interconnect_0_clock_crossing_io_s0_writedata),          //                                                   .writedata
		.clock_crossing_io_s0_burstcount                          (mm_interconnect_0_clock_crossing_io_s0_burstcount),         //                                                   .burstcount
		.clock_crossing_io_s0_byteenable                          (mm_interconnect_0_clock_crossing_io_s0_byteenable),         //                                                   .byteenable
		.clock_crossing_io_s0_readdatavalid                       (mm_interconnect_0_clock_crossing_io_s0_readdatavalid),      //                                                   .readdatavalid
		.clock_crossing_io_s0_waitrequest                         (mm_interconnect_0_clock_crossing_io_s0_waitrequest),        //                                                   .waitrequest
		.clock_crossing_io_s0_debugaccess                         (mm_interconnect_0_clock_crossing_io_s0_debugaccess),        //                                                   .debugaccess
		.cpu_jtag_debug_module_address                            (mm_interconnect_0_cpu_jtag_debug_module_address),           //                              cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                              (mm_interconnect_0_cpu_jtag_debug_module_write),             //                                                   .write
		.cpu_jtag_debug_module_read                               (mm_interconnect_0_cpu_jtag_debug_module_read),              //                                                   .read
		.cpu_jtag_debug_module_readdata                           (mm_interconnect_0_cpu_jtag_debug_module_readdata),          //                                                   .readdata
		.cpu_jtag_debug_module_writedata                          (mm_interconnect_0_cpu_jtag_debug_module_writedata),         //                                                   .writedata
		.cpu_jtag_debug_module_byteenable                         (mm_interconnect_0_cpu_jtag_debug_module_byteenable),        //                                                   .byteenable
		.cpu_jtag_debug_module_waitrequest                        (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),       //                                                   .waitrequest
		.cpu_jtag_debug_module_debugaccess                        (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),       //                                                   .debugaccess
		.jtag_uart_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                   .write
		.jtag_uart_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                   .read
		.jtag_uart_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                   .chipselect
		.onchip_memory2_s1_address                                (mm_interconnect_0_onchip_memory2_s1_address),               //                                  onchip_memory2_s1.address
		.onchip_memory2_s1_write                                  (mm_interconnect_0_onchip_memory2_s1_write),                 //                                                   .write
		.onchip_memory2_s1_readdata                               (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                                   .readdata
		.onchip_memory2_s1_writedata                              (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                                   .writedata
		.onchip_memory2_s1_byteenable                             (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                                   .byteenable
		.onchip_memory2_s1_chipselect                             (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                                   .chipselect
		.onchip_memory2_s1_clken                                  (mm_interconnect_0_onchip_memory2_s1_clken),                 //                                                   .clken
		.sma_in_s1_address                                        (mm_interconnect_0_sma_in_s1_address),                       //                                          sma_in_s1.address
		.sma_in_s1_readdata                                       (mm_interconnect_0_sma_in_s1_readdata),                      //                                                   .readdata
		.sma_out_s1_address                                       (mm_interconnect_0_sma_out_s1_address),                      //                                         sma_out_s1.address
		.sma_out_s1_write                                         (mm_interconnect_0_sma_out_s1_write),                        //                                                   .write
		.sma_out_s1_readdata                                      (mm_interconnect_0_sma_out_s1_readdata),                     //                                                   .readdata
		.sma_out_s1_writedata                                     (mm_interconnect_0_sma_out_s1_writedata),                    //                                                   .writedata
		.sma_out_s1_chipselect                                    (mm_interconnect_0_sma_out_s1_chipselect)                    //                                                   .chipselect
	);

	DE2_115_SD_CARD_NIOS_mm_interconnect_1 mm_interconnect_1 (
		.altpll_c0_clk                                          (c0_out_clk_clk),                                    //                                        altpll_c0.clk
		.altpll_c2_clk                                          (c2_out_clk_clk),                                    //                                        altpll_c2.clk
		.clock_crossing_io_m0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                // clock_crossing_io_m0_reset_reset_bridge_in_reset.reset
		.epp_i2c_scl_reset_reset_bridge_in_reset_reset          (cpu_jtag_debug_module_reset_reset),                 //          epp_i2c_scl_reset_reset_bridge_in_reset.reset
		.ir_reset_reset_bridge_in_reset_reset                   (rst_controller_003_reset_out_reset),                //                   ir_reset_reset_bridge_in_reset.reset
		.seg7_clock_sink_reset_reset_bridge_in_reset_reset      (rst_controller_001_reset_out_reset),                //      seg7_clock_sink_reset_reset_bridge_in_reset.reset
		.clock_crossing_io_m0_address                           (clock_crossing_io_m0_address),                      //                             clock_crossing_io_m0.address
		.clock_crossing_io_m0_waitrequest                       (clock_crossing_io_m0_waitrequest),                  //                                                 .waitrequest
		.clock_crossing_io_m0_burstcount                        (clock_crossing_io_m0_burstcount),                   //                                                 .burstcount
		.clock_crossing_io_m0_byteenable                        (clock_crossing_io_m0_byteenable),                   //                                                 .byteenable
		.clock_crossing_io_m0_read                              (clock_crossing_io_m0_read),                         //                                                 .read
		.clock_crossing_io_m0_readdata                          (clock_crossing_io_m0_readdata),                     //                                                 .readdata
		.clock_crossing_io_m0_readdatavalid                     (clock_crossing_io_m0_readdatavalid),                //                                                 .readdatavalid
		.clock_crossing_io_m0_write                             (clock_crossing_io_m0_write),                        //                                                 .write
		.clock_crossing_io_m0_writedata                         (clock_crossing_io_m0_writedata),                    //                                                 .writedata
		.clock_crossing_io_m0_debugaccess                       (clock_crossing_io_m0_debugaccess),                  //                                                 .debugaccess
		.epp_i2c_scl_s1_address                                 (mm_interconnect_1_epp_i2c_scl_s1_address),          //                                   epp_i2c_scl_s1.address
		.epp_i2c_scl_s1_write                                   (mm_interconnect_1_epp_i2c_scl_s1_write),            //                                                 .write
		.epp_i2c_scl_s1_readdata                                (mm_interconnect_1_epp_i2c_scl_s1_readdata),         //                                                 .readdata
		.epp_i2c_scl_s1_writedata                               (mm_interconnect_1_epp_i2c_scl_s1_writedata),        //                                                 .writedata
		.epp_i2c_scl_s1_chipselect                              (mm_interconnect_1_epp_i2c_scl_s1_chipselect),       //                                                 .chipselect
		.epp_i2c_sda_s1_address                                 (mm_interconnect_1_epp_i2c_sda_s1_address),          //                                   epp_i2c_sda_s1.address
		.epp_i2c_sda_s1_write                                   (mm_interconnect_1_epp_i2c_sda_s1_write),            //                                                 .write
		.epp_i2c_sda_s1_readdata                                (mm_interconnect_1_epp_i2c_sda_s1_readdata),         //                                                 .readdata
		.epp_i2c_sda_s1_writedata                               (mm_interconnect_1_epp_i2c_sda_s1_writedata),        //                                                 .writedata
		.epp_i2c_sda_s1_chipselect                              (mm_interconnect_1_epp_i2c_sda_s1_chipselect),       //                                                 .chipselect
		.i2c_scl_s1_address                                     (mm_interconnect_1_i2c_scl_s1_address),              //                                       i2c_scl_s1.address
		.i2c_scl_s1_write                                       (mm_interconnect_1_i2c_scl_s1_write),                //                                                 .write
		.i2c_scl_s1_readdata                                    (mm_interconnect_1_i2c_scl_s1_readdata),             //                                                 .readdata
		.i2c_scl_s1_writedata                                   (mm_interconnect_1_i2c_scl_s1_writedata),            //                                                 .writedata
		.i2c_scl_s1_chipselect                                  (mm_interconnect_1_i2c_scl_s1_chipselect),           //                                                 .chipselect
		.i2c_sda_s1_address                                     (mm_interconnect_1_i2c_sda_s1_address),              //                                       i2c_sda_s1.address
		.i2c_sda_s1_write                                       (mm_interconnect_1_i2c_sda_s1_write),                //                                                 .write
		.i2c_sda_s1_readdata                                    (mm_interconnect_1_i2c_sda_s1_readdata),             //                                                 .readdata
		.i2c_sda_s1_writedata                                   (mm_interconnect_1_i2c_sda_s1_writedata),            //                                                 .writedata
		.i2c_sda_s1_chipselect                                  (mm_interconnect_1_i2c_sda_s1_chipselect),           //                                                 .chipselect
		.ir_s1_address                                          (mm_interconnect_1_ir_s1_address),                   //                                            ir_s1.address
		.ir_s1_readdata                                         (mm_interconnect_1_ir_s1_readdata),                  //                                                 .readdata
		.key_s1_address                                         (mm_interconnect_1_key_s1_address),                  //                                           key_s1.address
		.key_s1_write                                           (mm_interconnect_1_key_s1_write),                    //                                                 .write
		.key_s1_readdata                                        (mm_interconnect_1_key_s1_readdata),                 //                                                 .readdata
		.key_s1_writedata                                       (mm_interconnect_1_key_s1_writedata),                //                                                 .writedata
		.key_s1_chipselect                                      (mm_interconnect_1_key_s1_chipselect),               //                                                 .chipselect
		.lcd_control_slave_address                              (mm_interconnect_1_lcd_control_slave_address),       //                                lcd_control_slave.address
		.lcd_control_slave_write                                (mm_interconnect_1_lcd_control_slave_write),         //                                                 .write
		.lcd_control_slave_read                                 (mm_interconnect_1_lcd_control_slave_read),          //                                                 .read
		.lcd_control_slave_readdata                             (mm_interconnect_1_lcd_control_slave_readdata),      //                                                 .readdata
		.lcd_control_slave_writedata                            (mm_interconnect_1_lcd_control_slave_writedata),     //                                                 .writedata
		.lcd_control_slave_begintransfer                        (mm_interconnect_1_lcd_control_slave_begintransfer), //                                                 .begintransfer
		.ledg_s1_address                                        (mm_interconnect_1_ledg_s1_address),                 //                                          ledg_s1.address
		.ledg_s1_write                                          (mm_interconnect_1_ledg_s1_write),                   //                                                 .write
		.ledg_s1_readdata                                       (mm_interconnect_1_ledg_s1_readdata),                //                                                 .readdata
		.ledg_s1_writedata                                      (mm_interconnect_1_ledg_s1_writedata),               //                                                 .writedata
		.ledg_s1_chipselect                                     (mm_interconnect_1_ledg_s1_chipselect),              //                                                 .chipselect
		.ledr_s1_address                                        (mm_interconnect_1_ledr_s1_address),                 //                                          ledr_s1.address
		.ledr_s1_write                                          (mm_interconnect_1_ledr_s1_write),                   //                                                 .write
		.ledr_s1_readdata                                       (mm_interconnect_1_ledr_s1_readdata),                //                                                 .readdata
		.ledr_s1_writedata                                      (mm_interconnect_1_ledr_s1_writedata),               //                                                 .writedata
		.ledr_s1_chipselect                                     (mm_interconnect_1_ledr_s1_chipselect),              //                                                 .chipselect
		.rs232_s1_address                                       (mm_interconnect_1_rs232_s1_address),                //                                         rs232_s1.address
		.rs232_s1_write                                         (mm_interconnect_1_rs232_s1_write),                  //                                                 .write
		.rs232_s1_read                                          (mm_interconnect_1_rs232_s1_read),                   //                                                 .read
		.rs232_s1_readdata                                      (mm_interconnect_1_rs232_s1_readdata),               //                                                 .readdata
		.rs232_s1_writedata                                     (mm_interconnect_1_rs232_s1_writedata),              //                                                 .writedata
		.rs232_s1_begintransfer                                 (mm_interconnect_1_rs232_s1_begintransfer),          //                                                 .begintransfer
		.rs232_s1_chipselect                                    (mm_interconnect_1_rs232_s1_chipselect),             //                                                 .chipselect
		.sd_clk_s1_address                                      (mm_interconnect_1_sd_clk_s1_address),               //                                        sd_clk_s1.address
		.sd_clk_s1_write                                        (mm_interconnect_1_sd_clk_s1_write),                 //                                                 .write
		.sd_clk_s1_readdata                                     (mm_interconnect_1_sd_clk_s1_readdata),              //                                                 .readdata
		.sd_clk_s1_writedata                                    (mm_interconnect_1_sd_clk_s1_writedata),             //                                                 .writedata
		.sd_clk_s1_chipselect                                   (mm_interconnect_1_sd_clk_s1_chipselect),            //                                                 .chipselect
		.sd_cmd_s1_address                                      (mm_interconnect_1_sd_cmd_s1_address),               //                                        sd_cmd_s1.address
		.sd_cmd_s1_write                                        (mm_interconnect_1_sd_cmd_s1_write),                 //                                                 .write
		.sd_cmd_s1_readdata                                     (mm_interconnect_1_sd_cmd_s1_readdata),              //                                                 .readdata
		.sd_cmd_s1_writedata                                    (mm_interconnect_1_sd_cmd_s1_writedata),             //                                                 .writedata
		.sd_cmd_s1_chipselect                                   (mm_interconnect_1_sd_cmd_s1_chipselect),            //                                                 .chipselect
		.sd_dat_s1_address                                      (mm_interconnect_1_sd_dat_s1_address),               //                                        sd_dat_s1.address
		.sd_dat_s1_write                                        (mm_interconnect_1_sd_dat_s1_write),                 //                                                 .write
		.sd_dat_s1_readdata                                     (mm_interconnect_1_sd_dat_s1_readdata),              //                                                 .readdata
		.sd_dat_s1_writedata                                    (mm_interconnect_1_sd_dat_s1_writedata),             //                                                 .writedata
		.sd_dat_s1_chipselect                                   (mm_interconnect_1_sd_dat_s1_chipselect),            //                                                 .chipselect
		.sd_wp_n_s1_address                                     (mm_interconnect_1_sd_wp_n_s1_address),              //                                       sd_wp_n_s1.address
		.sd_wp_n_s1_readdata                                    (mm_interconnect_1_sd_wp_n_s1_readdata),             //                                                 .readdata
		.seg7_avalon_slave_address                              (mm_interconnect_1_seg7_avalon_slave_address),       //                                seg7_avalon_slave.address
		.seg7_avalon_slave_write                                (mm_interconnect_1_seg7_avalon_slave_write),         //                                                 .write
		.seg7_avalon_slave_read                                 (mm_interconnect_1_seg7_avalon_slave_read),          //                                                 .read
		.seg7_avalon_slave_readdata                             (mm_interconnect_1_seg7_avalon_slave_readdata),      //                                                 .readdata
		.seg7_avalon_slave_writedata                            (mm_interconnect_1_seg7_avalon_slave_writedata),     //                                                 .writedata
		.sw_s1_address                                          (mm_interconnect_1_sw_s1_address),                   //                                            sw_s1.address
		.sw_s1_write                                            (mm_interconnect_1_sw_s1_write),                     //                                                 .write
		.sw_s1_readdata                                         (mm_interconnect_1_sw_s1_readdata),                  //                                                 .readdata
		.sw_s1_writedata                                        (mm_interconnect_1_sw_s1_writedata),                 //                                                 .writedata
		.sw_s1_chipselect                                       (mm_interconnect_1_sw_s1_chipselect),                //                                                 .chipselect
		.timer_s1_address                                       (mm_interconnect_1_timer_s1_address),                //                                         timer_s1.address
		.timer_s1_write                                         (mm_interconnect_1_timer_s1_write),                  //                                                 .write
		.timer_s1_readdata                                      (mm_interconnect_1_timer_s1_readdata),               //                                                 .readdata
		.timer_s1_writedata                                     (mm_interconnect_1_timer_s1_writedata),              //                                                 .writedata
		.timer_s1_chipselect                                    (mm_interconnect_1_timer_s1_chipselect),             //                                                 .chipselect
		.to_hw_port_s1_address                                  (mm_interconnect_1_to_hw_port_s1_address),           //                                    to_hw_port_s1.address
		.to_hw_port_s1_write                                    (mm_interconnect_1_to_hw_port_s1_write),             //                                                 .write
		.to_hw_port_s1_readdata                                 (mm_interconnect_1_to_hw_port_s1_readdata),          //                                                 .readdata
		.to_hw_port_s1_writedata                                (mm_interconnect_1_to_hw_port_s1_writedata),         //                                                 .writedata
		.to_hw_port_s1_chipselect                               (mm_interconnect_1_to_hw_port_s1_chipselect),        //                                                 .chipselect
		.to_hw_sig_s1_address                                   (mm_interconnect_1_to_hw_sig_s1_address),            //                                     to_hw_sig_s1.address
		.to_hw_sig_s1_write                                     (mm_interconnect_1_to_hw_sig_s1_write),              //                                                 .write
		.to_hw_sig_s1_readdata                                  (mm_interconnect_1_to_hw_sig_s1_readdata),           //                                                 .readdata
		.to_hw_sig_s1_writedata                                 (mm_interconnect_1_to_hw_sig_s1_writedata),          //                                                 .writedata
		.to_hw_sig_s1_chipselect                                (mm_interconnect_1_to_hw_sig_s1_chipselect),         //                                                 .chipselect
		.to_sw_sig_s1_address                                   (mm_interconnect_1_to_sw_sig_s1_address),            //                                     to_sw_sig_s1.address
		.to_sw_sig_s1_readdata                                  (mm_interconnect_1_to_sw_sig_s1_readdata)            //                                                 .readdata
	);

	DE2_115_SD_CARD_NIOS_irq_mapper irq_mapper (
		.clk           (c0_out_clk_clk),                     //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                    // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_50_clk_in_clk),                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_req      (),                                  // (terminated)
		.reset_req_in0  (1'b0),                              // (terminated)
		.reset_req_in1  (1'b0),                              // (terminated)
		.reset_in2      (1'b0),                              // (terminated)
		.reset_req_in2  (1'b0),                              // (terminated)
		.reset_in3      (1'b0),                              // (terminated)
		.reset_req_in3  (1'b0),                              // (terminated)
		.reset_in4      (1'b0),                              // (terminated)
		.reset_req_in4  (1'b0),                              // (terminated)
		.reset_in5      (1'b0),                              // (terminated)
		.reset_req_in5  (1'b0),                              // (terminated)
		.reset_in6      (1'b0),                              // (terminated)
		.reset_req_in6  (1'b0),                              // (terminated)
		.reset_in7      (1'b0),                              // (terminated)
		.reset_req_in7  (1'b0),                              // (terminated)
		.reset_in8      (1'b0),                              // (terminated)
		.reset_req_in8  (1'b0),                              // (terminated)
		.reset_in9      (1'b0),                              // (terminated)
		.reset_req_in9  (1'b0),                              // (terminated)
		.reset_in10     (1'b0),                              // (terminated)
		.reset_req_in10 (1'b0),                              // (terminated)
		.reset_in11     (1'b0),                              // (terminated)
		.reset_req_in11 (1'b0),                              // (terminated)
		.reset_in12     (1'b0),                              // (terminated)
		.reset_req_in12 (1'b0),                              // (terminated)
		.reset_in13     (1'b0),                              // (terminated)
		.reset_req_in13 (1'b0),                              // (terminated)
		.reset_in14     (1'b0),                              // (terminated)
		.reset_req_in14 (1'b0),                              // (terminated)
		.reset_in15     (1'b0),                              // (terminated)
		.reset_req_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk            (c0_out_clk_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (c2_out_clk_clk),                     //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (c0_out_clk_clk),                         //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_003_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
